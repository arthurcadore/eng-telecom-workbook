library ieee