s1 std_logic_vector(8 downto 0)

s1 <= std_logic_vector(to_unsigned(255,9))

